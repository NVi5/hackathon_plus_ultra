
module vio (
	source,
	probe);	

	output	[0:0]	source;
	input	[7:0]	probe;
endmodule
